module gpr (
				input clk, 
            input write_enable,
            input [4:0] AddrA,
            input [4:0] AddrB,
            input [4:0] AddrC, 
            output [31:0] A_out,        
            output [31:0] B_out,    
            input [31:0] C_in 
); 
// input and output initialization


reg [31:0] gpr [0:31]; // register array creation

initial begin
        $readmemb("values.txt", gpr); //reading from the file
end


always @(posedge clk) // posedge for clock value
begin
   gpr[5'b00000] <= 0; // $0 becomes 0 always 
   if(write_enable && AddrC != 0) 
        begin
            gpr[AddrC] <= C_in; 
        end
end

assign A_out = gpr[AddrA]; 
assign B_out = gpr[AddrB];

endmodule





////////////////////////

module testbench();

reg clk = 0;
reg write_enable = 1;
reg [4:0]AddrA;
reg [4:0]AddrB;
reg [4:0]AddrC;
reg [31:0] C_in;
wire [31:0]A_out;
wire [31:0]B_out;

gpr gpr (.clk(clk), .AddrA(AddrA), .AddrB(AddrB), 
			.AddrC(AddrC), .C_in(C_in), .A_out(A_out), .B_out(B_out),
			.write_enable(write_enable));

always begin 
#5;    clk = ~clk;
    
end
     
initial begin     
     AddrA = 5'b00000;
     AddrB = 5'b00010;
     AddrC = 5'b00110;
     C_in = 32'b00010_01100_10010_00000_10000_00000_01;


     #10;
     

     AddrA = 5'b01001;
     AddrB = 5'b10010;
     AddrC = 5'b01001;
     C_in = 32'b00010_01100_11110_00000_10000_00111_11;

     #10;
     

	  AddrA = 5'b11100;
     AddrB = 5'b00110;
     AddrC = 5'b01010;
     C_in = 32'b00010_00000_10010_00000_10000_00000_01;

     #10;
     

     AddrA = 5'b01001;
     AddrB = 5'b11111;
     AddrC = 5'b01001;
     C_in = 32'b00010_01100_11110_11111_10000_00111_11;

     #10;
end
     
endmodule




///////////_Values.txt_////////
00000000000000001111111100000000
00000000000000000000000000000000
00000000000001010101010100000000
00000000000000001000000000000000
00000000000000000000010000000000
00011111100000000000000000000000
00000000000000111100000000000000
00000001010000000000000000000000
00000000000001010101001100000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000001010101001100000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000001010101001100000000
00000000000000000000000000000000
00011111100000000000000000000000
00000000000001010101001100000000
00011111100000000000000000000000
00000000000001010101001100000000
00000000000001010101001100000000
00000000000000001111111100000000
00000000000001010101010100000000
00000000000000000000000000000000
00000000000000000000000000000000
00111110000000000000001111111000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000001010101010100000000


